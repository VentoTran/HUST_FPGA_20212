LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

ENTITY TEST_KIT IS
	PORT(
		CLK				: IN		STD_LOGIC;
		SW					: IN		STD_LOGIC_VECTOR (9 DOWNTO 0);
		LEDR				: OUT		STD_LOGIC_VECTOR (9 DOWNTO 0);
		KEY				: IN		STD_LOGIC_VECTOR (3 DOWNTO 0);
		LEDG				: OUT 	STD_LOGIC_VECTOR (7 DOWNTO 0);
		LED7_0			: OUT		STD_LOGIC_VECTOR (6 DOWNTO 0);
		LED7_1			: OUT		STD_LOGIC_VECTOR (6 DOWNTO 0);
		LED7_2			: OUT		STD_LOGIC_VECTOR (6 DOWNTO 0);
		LED7_3			: OUT		STD_LOGIC_VECTOR (6 DOWNTO 0)
	);
END TEST_KIT;



ARCHITECTURE BEHAVIOUR OF TEST_KIT IS

	SIGNAL i	:	INTEGER RANGE 0 TO 15;
	
	TYPE ARR6bLED7A IS ARRAY (1 to 10) OF STD_LOGIC_VECTOR(6 DOWNTO 0);
	CONSTANT LED7A	:	ARR6bLED7A	:=	("1000000","1111001","0100100","0110000","0011001","0010010","0000010","1111000","0000000","0010000");
	
BEGIN

	PROCESS (CLK)
	BEGIN
		IF (CLK'EVENT AND CLK = '1') THEN
		
			LEDR <= SW;
			i <= 15 - to_integer(unsigned(KEY));
			LEDG <= std_logic_vector(to_unsigned(i, LEDG'length));
			IF (i < 10) THEN
				LED7_0 <= LED7A(i+1)(6 DOWNTO 0);
			END IF;
		
		END IF;
	END PROCESS;



END BEHAVIOUR;